library ieee;
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;

entity ROM_176x4 is
  port (Clock : in std_logic;
  		CS_L : in std_logic;
        R_W  : in std_logic;
        Addr   : in std_logic_vector(7 downto 0);
        Data  : out std_logic_vector(3 downto 0));
end ROM_176x4;

architecture ROM_176x4_Arch of ROM_176x4 is
  type rom_type is array (0 to 175)
        of std_logic_vector (3 downto 0);
  signal ROM : rom_type;
  signal Read_Enable : std_logic;
begin

ROM(0) <= X"7";
ROM(1) <= X"0";
ROM(2) <= X"D";
ROM(3) <= X"0";
ROM(4) <= X"B";
ROM(5) <= X"D";
ROM(6) <= X"1";
ROM(7) <= X"B";
ROM(8) <= X"5";
ROM(9) <= X"0";
ROM(10) <= X"B";
ROM(11) <= X"5";
ROM(12) <= X"2";
ROM(13) <= X"9";
ROM(14) <= X"0";
ROM(15) <= X"1";
ROM(16) <= X"F";
ROM(17) <= X"0";
ROM(18) <= X"B";
ROM(19) <= X"6";
ROM(20) <= X"1";
ROM(21) <= X"D";
ROM(22) <= X"0";
ROM(23) <= X"B";
ROM(24) <= X"6";
ROM(25) <= X"6";
ROM(26) <= X"A";
ROM(27) <= X"E";
ROM(28) <= X"3";
ROM(29) <= X"F";
ROM(30) <= X"0";
ROM(31) <= X"B";
ROM(32) <= X"4";
ROM(33) <= X"2";
ROM(34) <= X"9";
ROM(35) <= X"8";
ROM(36) <= X"0";
ROM(37) <= X"7";
ROM(38) <= X"1";
ROM(39) <= X"1";
ROM(40) <= X"E";
ROM(41) <= X"0";
ROM(42) <= X"B";
ROM(43) <= X"D";
ROM(44) <= X"0";
ROM(45) <= X"B";
ROM(46) <= X"6";
ROM(47) <= X"1";
ROM(48) <= X"A";
ROM(49) <= X"7";
ROM(50) <= X"6";
ROM(51) <= X"F";
ROM(52) <= X"0";
ROM(53) <= X"B";
ROM(54) <= X"4";
ROM(55) <= X"2";
ROM(56) <= X"A";
ROM(57) <= X"7";
ROM(58) <= X"6";
ROM(59) <= X"9";
ROM(60) <= X"8";
ROM(61) <= X"0";
ROM(62) <= X"F";
ROM(63) <= X"1";
ROM(64) <= X"B";
ROM(65) <= X"6";
ROM(66) <= X"1";
ROM(67) <= X"D";
ROM(68) <= X"1";
ROM(69) <= X"B";
ROM(70) <= X"7";
ROM(71) <= X"0";
ROM(72) <= X"D";
ROM(73) <= X"0";
ROM(74) <= X"B";
ROM(75) <= X"4";
ROM(76) <= X"2";
ROM(77) <= X"F";
ROM(78) <= X"1";
ROM(79) <= X"B";
ROM(80) <= X"6";
ROM(81) <= X"6";
ROM(82) <= X"A";
ROM(83) <= X"D";
ROM(84) <= X"5";
ROM(85) <= X"F";
ROM(86) <= X"1";
ROM(87) <= X"B";
ROM(88) <= X"4";
ROM(89) <= X"1";
ROM(90) <= X"9";
ROM(91) <= X"8";
ROM(92) <= X"0";
ROM(93) <= X"7";
ROM(94) <= X"0";
ROM(95) <= X"D";
ROM(96) <= X"1";
ROM(97) <= X"B";
ROM(98) <= X"4";
ROM(99) <= X"1";
ROM(100) <= X"9";
ROM(101) <= X"8";
ROM(102) <= X"0";
ROM(103) <= X"7";
ROM(104) <= X"9";
ROM(105) <= X"D";
ROM(106) <= X"0";
ROM(107) <= X"B";
ROM(108) <= X"4";
ROM(109) <= X"2";
ROM(110) <= X"7";
ROM(111) <= X"1";
ROM(112) <= X"1";
ROM(113) <= X"E";
ROM(114) <= X"1";
ROM(115) <= X"B";
ROM(116) <= X"6";
ROM(117) <= X"1";
ROM(118) <= X"A";
ROM(119) <= X"E";
ROM(120) <= X"7";
ROM(121) <= X"F";
ROM(122) <= X"1";
ROM(123) <= X"B";
ROM(124) <= X"4";
ROM(125) <= X"1";
ROM(126) <= X"7";
ROM(127) <= X"9";
ROM(128) <= X"D";
ROM(129) <= X"1";
ROM(130) <= X"B";
ROM(131) <= X"4";
ROM(132) <= X"1";
ROM(133) <= X"9";
ROM(134) <= X"8";
ROM(135) <= X"0";
ROM(136) <= X"0";
ROM(137) <= X"0";
ROM(138) <= X"0";
ROM(139) <= X"0";
ROM(140) <= X"0";
ROM(141) <= X"0";
ROM(142) <= X"0";
ROM(143) <= X"0";
ROM(144) <= X"0";
ROM(145) <= X"0";
ROM(146) <= X"0";
ROM(147) <= X"0";
ROM(148) <= X"0";
ROM(149) <= X"0";
ROM(150) <= X"0";
ROM(151) <= X"0";
ROM(152) <= X"0";
ROM(153) <= X"0";
ROM(154) <= X"0";
ROM(155) <= X"0";
ROM(156) <= X"0";
ROM(157) <= X"0";
ROM(158) <= X"0";
ROM(159) <= X"0";
ROM(160) <= X"0";
ROM(161) <= X"0";
ROM(162) <= X"0";
ROM(163) <= X"0";
ROM(164) <= X"0";
ROM(165) <= X"0";
ROM(166) <= X"0";
ROM(167) <= X"0";
ROM(168) <= X"0";
ROM(169) <= X"0";
ROM(170) <= X"0";
ROM(171) <= X"0";
ROM(172) <= X"0";
ROM(173) <= X"0";
ROM(174) <= X"0";
ROM(175) <= X"0";
	Read_Enable <=  '0' when(CS_L='0' and R_W = '1') else '1';

	process (Clock)
	begin
		if(Clock='0') then
			if(Read_Enable = '0') then
			  Data  <= ROM(conv_integer(Addr));
		  	else
			  Data <= "ZZZZ";
	      	end if;
		else Data <= "ZZZZ";
		end if;

	end process;

	end ROM_176x4_Arch;
